// ECE:3350 SISC processor project
// main SISC module, part 1
// Nick Smith and Alan Rolla

`timescale 1ns/100ps  

module sisc (clk, rst_f, ir);

  input clk, rst_f;
  input [31:0] ir;

// declare all internal wires here
	wire [1:0] ALU_OP;
	wire WB_SEL;
	wire RF_WE;
	wire STAT_EN;
	wire 

// component instantiation goes here


  initial
  
// put a $monitor statement here.  



endmodule


